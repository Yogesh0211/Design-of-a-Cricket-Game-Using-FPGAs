module cricketGame(
    input clk_fpga,
    input reset,
    input delivery,
    input teamSwitch,
    output [7:0] runs,
    output [3:0] wickets,
    output [7:0] leds,
    output inningOver,
    output gameOver,
    output winner
    );
	 
	 wire [11:0] team1Data; // stores and updates teaml's runs and wickets when switch is 0 
	 wire [11:0] team2Data; // stores and updates team2's runs and wickets when switch is 1 
	 wire [6:0] team1Balls; // the number of teaml's deliveries that are legal balls, shown on LEDs 
	 wire [6:0] team2Balls; // the number of team2's deliveries that are legal balls, shown on LEDs 
	 wire [3:0] lfsr_out;   // pseudorandom number from linear feedback shift register
	 
	 // pseudo random number generator using a linear feedback shift register 
	 lfsr g1(clk_fgpa, reset, lfsr_out);
	 // assign score and wickets based on pseudo random number generated by lfsr 
	 score_and_wickets g2(clk_fpga, reset, delivery, teamSwitch, lfsr_out, gameOver, runs, wickets, team1Data, team2Data);
	 // comparator that finds and locks in the winner when the game is over 
	 score_comparator g3(clk_fpga, reset, team1Data, team2Data, team1Balls, team2Balls, wickets, leds, inningOver, gameOver, winner);
	 // assign Leds based on balls of team in play, or scroll leds when the game is over 
	 led_controller g4(clk_fpga, reset, teamSwitch, delivery, lfsr_out, inningOver, gameOver, leds, team1Balls, team2Balls);

endmodule
